/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_WillyJules_chipbootcamp (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

assign uio_out = 0;
  assign uio_oe  = 0;

  // Coordinates
  reg [3:0] x0, y0, x1, y1;
  reg [3:0] x, y;
  reg [4:0] dx, dy, err, sx, sy; // 5 bits to prevent overflow
  reg done;

  always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      x0 <= ui_in[7:4];
      y0 <= ui_in[3:0];
      x1 <= uio_in[7:4];
      y1 <= uio_in[3:0];

      x <= ui_in[7:4];
      y <= ui_in[3:0];

      dx <= (uio_in[7:4] > ui_in[7:4]) ? (uio_in[7:4] - ui_in[7:4]) : (ui_in[7:4] - uio_in[7:4]);
      dy <= (uio_in[3:0] > ui_in[3:0]) ? (uio_in[3:0] - ui_in[3:0]) : (ui_in[3:0] - uio_in[3:0]);
      
      sx <= (ui_in[7:4] < uio_in[7:4]) ? 1 : -1;
      sy <= (ui_in[3:0] < uio_in[3:0]) ? 1 : -1;

      err <= (dx > dy) ? (dx >> 1) : -(dy >> 1);
      done <= 0;
    end else if (!done) begin
      // Output current coordinate
      uo_out <= {x, y};

      if ((x == x1) && (y == y1)) begin
        done <= 1;
      end else begin
        reg [4:0] e2;
        e2 = err;
        if (e2 > -dx) begin
          err <= err - dy;
          x <= x + sx[0]; // convert sx to 0/1
        end
        if (e2 < dy) begin
          err <= err + dx;
          y <= y + sy[0];
        end
      end
    end
  end
  // List all unused inputs to prevent warnings
  wire _unused = &{ena, clk, rst_n, 1'b0};

endmodule
